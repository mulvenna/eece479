magic
tech scmos
timestamp 1428795988
<< pwell >>
rect 4098 361 4144 377
rect 4048 341 4084 355
rect 4009 221 4043 233
<< nwell >>
rect 4098 384 4146 395
rect 4049 359 4085 373
rect 4010 246 4044 258
<< polysilicon >>
rect -22 781 6 783
rect 2614 781 2698 783
rect -22 82 -18 781
rect 2398 717 2403 719
rect 95 647 2417 649
rect 4116 390 4119 392
rect 4116 373 4119 387
rect 4066 366 4069 369
rect 4116 368 4119 370
rect 4066 359 4069 363
rect 4066 355 4068 359
rect 4066 351 4069 355
rect 4066 345 4069 348
rect 3990 297 4024 300
rect 3990 288 4003 291
rect 4000 254 4003 288
rect 4022 252 4024 297
rect 4022 242 4024 248
rect 4022 239 4070 242
rect 4022 231 4024 239
rect 4022 225 4024 227
rect 2611 82 2614 99
rect -22 79 6 82
<< ndiffusion >>
rect 4114 370 4116 373
rect 4119 370 4121 373
rect 4063 348 4066 351
rect 4069 348 4073 351
rect 4020 227 4022 231
rect 4024 227 4026 231
<< pdiffusion >>
rect 4114 387 4116 390
rect 4119 387 4121 390
rect 4063 363 4066 366
rect 4069 363 4072 366
rect 4020 248 4022 252
rect 4024 248 4026 252
<< metal1 >>
rect 83 862 92 865
rect 392 862 417 865
rect 719 862 744 865
rect 1043 862 1070 865
rect 1370 862 1395 865
rect 1696 862 1721 865
rect 2022 862 2047 865
rect 2348 862 2373 865
rect 83 838 86 862
rect 2543 839 2555 843
rect 2582 826 2615 829
rect 2582 793 2585 826
rect 2664 810 2677 814
rect 2663 801 2673 805
rect 2544 789 2567 792
rect 2605 786 2614 790
rect 2679 790 2698 794
rect 172 618 2643 622
rect 2639 545 2643 618
rect 2743 545 2749 548
rect 2639 541 2749 545
rect 2684 403 2688 419
rect 2698 417 2702 419
rect 2698 403 2702 413
rect 2712 403 2716 415
rect 2856 403 2860 419
rect 2870 417 2874 419
rect 2870 403 2874 413
rect 2884 403 2888 415
rect 3028 403 3032 419
rect 3042 417 3046 419
rect 3042 403 3046 413
rect 3056 403 3060 415
rect 3200 403 3204 419
rect 3214 417 3218 419
rect 3214 403 3218 413
rect 3228 403 3232 415
rect 3372 403 3376 419
rect 3386 417 3390 419
rect 3386 403 3390 413
rect 3400 403 3404 415
rect 3544 403 3548 419
rect 3558 417 3562 419
rect 3558 403 3562 413
rect 3572 403 3576 415
rect 3716 403 3720 412
rect 3730 403 3734 413
rect 3744 403 3748 415
rect 3888 403 3892 417
rect 3902 403 3906 413
rect 3916 403 3920 415
rect 3990 396 4164 400
rect 3990 387 4079 391
rect 4075 383 4079 387
rect 4125 387 4130 391
rect 4134 388 4139 391
rect 4110 383 4114 387
rect 3990 380 3997 381
rect 4075 380 4114 383
rect 3990 377 4066 380
rect 4062 376 4066 377
rect 4062 373 4104 376
rect 3990 367 4055 371
rect 3990 357 4036 361
rect 3935 330 4015 334
rect 4031 329 4036 357
rect 4051 359 4055 367
rect 4076 364 4080 367
rect 4084 364 4090 367
rect 4059 359 4063 363
rect 4051 356 4063 359
rect 4059 352 4063 356
rect 4072 356 4084 359
rect 4073 344 4076 348
rect 4073 336 4076 340
rect 4081 329 4084 356
rect 4100 346 4104 373
rect 4110 374 4114 380
rect 4123 379 4153 383
rect 4121 366 4125 370
rect 3989 313 3995 327
rect 4031 326 4111 329
rect 4121 321 4125 362
rect 4137 326 4148 330
rect 4077 317 4125 321
rect 3989 309 4148 313
rect 3990 262 4072 266
rect 4027 259 4030 262
rect 4027 255 4036 259
rect 2567 245 2571 249
rect 2558 242 2571 245
rect 4027 252 4030 255
rect 4000 242 4004 250
rect 4016 242 4020 248
rect 4000 239 4020 242
rect 4016 231 4020 239
rect 4026 225 4030 227
rect 4026 222 4036 225
rect 4040 222 4052 226
rect 4026 221 4030 222
rect 175 41 179 57
rect 501 41 505 57
rect 827 40 831 56
rect 1153 41 1157 57
rect 1479 38 1483 54
rect 1805 39 1809 55
rect 2131 40 2135 56
rect 2457 39 2462 49
rect 2706 41 2710 57
rect 2878 42 2882 58
rect 3050 41 3054 57
rect 3222 40 3226 56
rect 3394 48 3398 56
rect 3566 40 3570 56
rect 3738 48 3742 56
rect 3910 48 3914 56
<< metal2 >>
rect 2553 835 2605 839
rect 2571 789 2581 793
rect 2601 790 2605 835
rect 2674 794 2679 800
rect 121 745 339 749
rect 447 745 665 749
rect 773 745 991 749
rect 1099 745 1317 749
rect 1425 745 1643 749
rect 1751 745 1969 749
rect 2077 745 2295 749
rect 2674 592 2679 789
rect 2553 589 2679 592
rect 2553 259 2558 589
rect 2712 471 3990 475
rect 2712 419 2716 471
rect 2688 413 2698 417
rect 2884 463 3990 467
rect 2884 419 2888 463
rect 2860 413 2870 417
rect 3056 455 3990 459
rect 3056 419 3060 455
rect 3032 413 3042 417
rect 3228 447 3990 451
rect 3228 419 3232 447
rect 3204 413 3214 417
rect 3400 439 3990 443
rect 3400 419 3404 439
rect 3376 413 3386 417
rect 3572 431 3990 435
rect 3572 419 3576 431
rect 3548 413 3558 417
rect 3744 423 3990 427
rect 3744 419 3748 423
rect 3720 413 3730 417
rect 3892 414 3902 417
rect 3920 415 3990 419
rect 4090 354 4094 364
rect 4130 354 4134 387
rect 4090 351 4134 354
rect 4015 327 4019 330
rect 4073 327 4076 332
rect 4015 324 4076 327
rect 4073 321 4076 324
rect 4073 298 4077 317
rect 4052 295 4077 298
rect 2553 245 2557 259
rect 4052 226 4056 295
rect 4090 265 4094 351
rect 4139 346 4142 375
rect 4104 342 4142 346
rect 4115 326 4133 330
rect 4076 262 4094 265
<< ntransistor >>
rect 4116 370 4119 373
rect 4066 348 4069 351
rect 4022 227 4024 231
<< ptransistor >>
rect 4116 387 4119 390
rect 4066 363 4069 366
rect 4022 248 4024 252
<< polycontact >>
rect 2610 806 2614 810
rect 292 770 296 774
rect 618 770 622 774
rect 944 770 948 774
rect 1270 770 1274 774
rect 1596 770 1600 774
rect 1922 770 1926 774
rect 2248 770 2252 774
rect 2574 769 2579 774
rect 4119 379 4123 383
rect 4068 355 4072 359
rect 2567 249 2571 253
rect 4000 250 4004 254
<< ndcontact >>
rect 4110 370 4114 374
rect 4121 370 4125 374
rect 4059 348 4063 352
rect 4073 348 4077 352
rect 4016 227 4020 231
rect 4026 227 4030 231
<< pdcontact >>
rect 4110 387 4114 391
rect 4121 387 4125 391
rect 4059 363 4063 367
rect 4072 363 4076 367
rect 4016 248 4020 252
rect 4026 248 4030 252
<< m2contact >>
rect 2673 800 2680 805
rect 2567 789 2571 793
rect 2581 789 2585 793
rect 2601 785 2605 790
rect 2674 789 2679 794
rect 167 618 172 622
rect 2698 413 2702 417
rect 2712 415 2716 419
rect 2870 413 2874 417
rect 2884 415 2888 419
rect 3042 413 3046 417
rect 3056 415 3060 419
rect 3214 413 3218 417
rect 3228 415 3232 419
rect 3386 413 3390 417
rect 3400 415 3404 419
rect 3558 413 3562 417
rect 3572 415 3576 419
rect 3730 413 3734 417
rect 3744 415 3748 419
rect 3902 413 3906 417
rect 3916 415 3920 419
rect 4130 387 4134 391
rect 4015 330 4019 334
rect 4090 364 4094 368
rect 4073 332 4077 336
rect 4139 375 4143 379
rect 4100 342 4104 346
rect 4111 326 4115 330
rect 4133 326 4137 330
rect 4073 317 4077 321
rect 4072 262 4076 266
rect 2553 241 2558 245
rect 4052 222 4056 226
<< psubstratepcontact >>
rect 4121 362 4125 366
rect 4073 340 4077 344
rect 4036 222 4040 226
<< nsubstratencontact >>
rect 4139 387 4143 391
rect 4080 364 4084 368
rect 4036 255 4040 259
use dbithigh  dbithigh_0
timestamp 1428795971
transform 1 0 100 0 1 796
box -94 -747 232 141
use dbithigh  dbithigh_1
timestamp 1428795971
transform 1 0 426 0 1 796
box -94 -747 232 141
use dbithigh  dbithigh_2
timestamp 1428795971
transform 1 0 752 0 1 796
box -94 -747 232 141
use dbithigh  dbithigh_3
timestamp 1428795971
transform 1 0 1078 0 1 796
box -94 -747 232 141
use dbithigh  dbithigh_4
timestamp 1428795971
transform 1 0 1404 0 1 796
box -94 -747 232 141
use dbithigh  dbithigh_5
timestamp 1428795971
transform 1 0 1730 0 1 796
box -94 -747 232 141
use dbithigh  dbithigh_6
timestamp 1428795971
transform 1 0 2056 0 1 796
box -94 -747 232 141
use dbithigh  dbithigh_7
timestamp 1428795971
transform 1 0 2382 0 1 796
box -94 -747 232 141
use ../cells/and  and_0
timestamp 1428029823
transform -1 0 2639 0 1 805
box -25 -19 25 24
use dbitlow  dbitlow_0
timestamp 1428705999
transform 1 0 2671 0 1 348
box -57 -292 116 69
use dbitlow  dbitlow_1
timestamp 1428705999
transform 1 0 2843 0 1 348
box -57 -292 116 69
use dbitlow  dbitlow_2
timestamp 1428705999
transform 1 0 3015 0 1 348
box -57 -292 116 69
use dbitlow  dbitlow_3
timestamp 1428705999
transform 1 0 3187 0 1 348
box -57 -292 116 69
use dbitlow  dbitlow_4
timestamp 1428705999
transform 1 0 3359 0 1 348
box -57 -292 116 69
use dbitlow  dbitlow_5
timestamp 1428705999
transform 1 0 3531 0 1 348
box -57 -292 116 69
use dbitlow  dbitlow_6
timestamp 1428705999
transform 1 0 3703 0 1 348
box -57 -292 116 69
use dbitlow  dbitlow_7
timestamp 1428705999
transform 1 0 3875 0 1 348
box -57 -292 116 69
<< labels >>
rlabel metal1 2675 812 2675 812 1 load
rlabel metal1 2672 803 2672 803 1 clk
rlabel metal1 4144 327 4144 327 1 sel2
rlabel metal1 4147 381 4147 381 1 sel1
rlabel polysilicon 121 648 121 648 1 add
rlabel metal1 4139 310 4139 310 1 inbit
rlabel metal1 4057 264 4057 264 1 Vdd
rlabel metal1 4061 399 4061 399 1 Gnd
rlabel polysilicon 4047 240 4047 240 1 shift
rlabel metal2 3987 473 3987 473 1 dividendin_7
rlabel metal2 3986 465 3986 465 1 dividendin_6
rlabel metal2 3985 457 3985 457 1 dividendin_5
rlabel metal2 3985 449 3985 449 1 dividendin_4
rlabel metal2 3985 441 3985 441 1 dividendin_3
rlabel metal2 3984 433 3984 433 1 dividendin_2
rlabel metal2 3983 426 3983 426 1 dividendin_1
rlabel metal2 3982 418 3982 418 1 dividendin_0
rlabel polysilicon -20 85 -20 85 3 reset
rlabel metal1 3912 51 3912 51 1 quotient_0
rlabel metal1 3739 51 3739 51 1 quotient_1
rlabel metal1 3567 49 3567 49 1 quotient_2
rlabel metal1 3396 51 3396 51 1 quotient_3
rlabel metal1 3223 51 3223 51 1 quotient_4
rlabel metal1 3051 50 3051 50 1 quotient_5
rlabel metal1 2881 51 2881 51 1 quotient_6
rlabel metal1 2707 51 2707 51 1 quotient_7
rlabel metal1 2133 44 2133 44 1 remainder_0
rlabel metal1 1806 44 1806 44 1 remainder_1
rlabel metal1 1481 42 1481 42 1 remainder_2
rlabel metal1 1154 45 1154 45 1 remainder_3
rlabel metal1 829 44 829 44 1 remainder_4
rlabel metal1 502 44 502 44 1 remainder_5
rlabel metal1 177 45 177 45 1 remainder_6
rlabel metal1 400 863 400 863 1 divisorin_6
rlabel metal1 726 863 726 863 1 divisorin_5
rlabel metal1 1056 864 1056 864 1 divisorin_4
rlabel metal1 1380 864 1380 864 1 divisorin_3
rlabel metal1 1706 864 1706 864 1 divisorin_2
rlabel metal1 2032 863 2032 863 1 divisorin_1
rlabel metal1 2359 864 2359 864 1 divisorin_0
rlabel metal1 2460 44 2460 44 1 hello
<< end >>
