magic
tech scmos
timestamp 1428726019
<< pwell >>
rect -13 0 64 17
<< nwell >>
rect -13 28 64 45
<< polysilicon >>
rect -4 38 -2 40
rect 5 38 7 40
rect 13 38 15 40
rect 21 38 23 40
rect 29 38 31 40
rect 54 38 56 40
rect -4 13 -2 32
rect 5 13 7 32
rect 13 13 15 32
rect 21 13 23 32
rect 29 13 31 32
rect 54 13 56 32
rect -4 8 -2 10
rect 5 8 7 10
rect 13 8 15 10
rect 21 8 23 10
rect 29 8 31 10
rect 54 8 56 10
<< ndiffusion >>
rect -6 10 -4 13
rect -2 10 5 13
rect 7 10 13 13
rect 15 10 21 13
rect 23 10 29 13
rect 31 10 33 13
rect 53 10 54 13
rect 56 10 58 13
<< pdiffusion >>
rect -6 32 -4 38
rect -2 32 0 38
rect 4 32 5 38
rect 7 32 8 38
rect 12 32 13 38
rect 15 32 16 38
rect 20 32 21 38
rect 23 32 24 38
rect 28 32 29 38
rect 31 32 33 38
rect 53 32 54 38
rect 56 32 58 38
<< metal1 >>
rect -10 42 9 44
rect 13 42 53 44
rect -10 41 53 42
rect -10 38 -6 41
rect 8 38 12 41
rect 24 38 28 41
rect 49 38 53 41
rect 0 25 4 32
rect 16 25 20 32
rect 33 25 37 32
rect 58 25 62 32
rect 0 22 50 25
rect 33 13 37 22
rect 58 22 66 25
rect 58 13 62 22
rect -10 6 -6 9
rect 49 6 53 9
rect -10 3 8 6
rect 12 3 53 6
<< ntransistor >>
rect -4 10 -2 13
rect 5 10 7 13
rect 13 10 15 13
rect 21 10 23 13
rect 29 10 31 13
rect 54 10 56 13
<< ptransistor >>
rect -4 32 -2 38
rect 5 32 7 38
rect 13 32 15 38
rect 21 32 23 38
rect 29 32 31 38
rect 54 32 56 38
<< polycontact >>
rect 50 21 54 25
<< ndcontact >>
rect -10 9 -6 13
rect 33 9 37 13
rect 49 9 53 13
rect 58 9 62 13
<< pdcontact >>
rect -10 32 -6 38
rect 0 32 4 38
rect 8 32 12 38
rect 16 32 20 38
rect 24 32 28 38
rect 33 32 37 38
rect 49 32 53 38
rect 58 32 62 38
<< psubstratepcontact >>
rect 8 2 12 6
<< nsubstratencontact >>
rect 9 42 13 46
<< labels >>
rlabel polysilicon -3 26 -3 26 1 a
rlabel polysilicon 6 20 6 20 1 b
rlabel polysilicon 14 20 14 20 1 c
rlabel polysilicon 22 20 22 20 1 d
rlabel polysilicon 30 20 30 20 1 e
rlabel metal1 19 4 19 4 1 Gnd
rlabel metal1 18 42 18 42 5 Vdd
rlabel metal1 64 23 64 23 7 q
<< end >>
