magic
tech scmos
timestamp 1428786523
<< pwell >>
rect -89 12 -49 25
rect 88 12 123 14
rect -89 4 123 12
rect -83 2 123 4
rect -83 -6 88 2
rect -113 -7 88 -6
rect -113 -23 145 -7
rect -48 -28 145 -23
rect -48 -31 88 -28
<< nwell >>
rect -48 53 88 61
rect -112 35 88 53
rect -112 33 146 35
rect -112 2 -93 33
rect -48 20 146 33
rect -48 18 88 20
rect 126 0 146 20
<< polysilicon >>
rect -35 50 -28 52
rect -24 50 11 52
rect 15 50 40 52
rect 43 50 74 52
rect 78 50 80 52
rect -82 40 -80 42
rect -82 21 -80 36
rect -82 15 -80 17
rect -82 13 -70 15
rect -57 13 -47 15
rect -72 9 -70 13
rect -102 7 -100 9
rect -72 7 -68 9
rect -102 2 -100 4
rect -102 0 -86 2
rect -102 -7 -100 0
rect -68 1 -66 5
rect -51 4 -47 13
rect -35 6 -33 50
rect 3 48 7 50
rect 65 48 69 50
rect -37 4 -33 6
rect -31 42 -28 44
rect -24 42 11 44
rect 15 42 49 44
rect 52 42 74 44
rect 78 42 80 44
rect -102 -12 -100 -10
rect -68 -15 -66 -2
rect -51 -9 -48 4
rect -37 -6 -35 4
rect -31 1 -29 42
rect 27 36 48 37
rect 27 35 58 36
rect 27 33 29 35
rect 46 34 58 35
rect 61 34 74 36
rect 78 34 80 36
rect -7 31 29 33
rect -7 29 -4 31
rect 29 26 34 28
rect 38 26 40 28
rect -7 8 -4 25
rect 29 17 31 26
rect 104 28 106 30
rect 104 23 106 25
rect 97 21 106 23
rect 26 15 31 17
rect 97 18 99 21
rect 94 16 99 18
rect -22 6 -4 8
rect -7 4 -4 6
rect 29 6 31 15
rect 104 13 106 21
rect 104 8 106 10
rect 29 4 34 6
rect 38 4 40 6
rect -7 -2 -4 0
rect -7 -3 25 -2
rect 91 -3 93 6
rect 133 5 135 7
rect 133 -3 135 2
rect -37 -8 -33 -6
rect -51 -15 -48 -12
rect -35 -20 -33 -8
rect -31 -12 -29 -3
rect -7 -4 60 -3
rect 23 -5 60 -4
rect 63 -5 74 -3
rect 23 -7 26 -5
rect 71 -6 74 -5
rect 78 -6 80 -3
rect 91 -5 135 -3
rect 133 -9 135 -5
rect -31 -14 -28 -12
rect -24 -14 11 -12
rect 15 -14 51 -12
rect 54 -14 74 -12
rect 78 -14 80 -12
rect 133 -14 135 -12
rect -35 -22 -28 -20
rect -24 -22 11 -20
rect 15 -22 40 -20
rect 43 -22 74 -20
rect 78 -22 80 -20
<< ndiffusion >>
rect -84 17 -82 21
rect -80 17 -77 21
rect -71 -2 -68 1
rect -66 -2 -60 1
rect -104 -10 -102 -7
rect -100 -10 -98 -7
rect 34 6 38 7
rect 103 10 104 13
rect 106 10 107 13
rect -8 0 -7 4
rect -4 0 -3 4
rect 34 3 38 4
rect 60 -3 63 -2
rect 74 -3 78 -2
rect -53 -12 -51 -9
rect -48 -12 -46 -9
rect -28 -12 -24 -11
rect 11 -12 15 -11
rect 51 -12 54 -10
rect 60 -7 63 -5
rect 74 -12 78 -6
rect 132 -12 133 -9
rect 135 -12 136 -9
rect -28 -15 -24 -14
rect -28 -20 -24 -19
rect 11 -20 15 -14
rect 51 -15 54 -14
rect 40 -20 43 -19
rect 74 -20 78 -14
rect -28 -23 -24 -22
rect 11 -23 15 -22
rect 40 -23 43 -22
rect 74 -23 78 -22
<< pdiffusion >>
rect -28 52 -24 53
rect 11 52 15 53
rect 40 52 43 53
rect 74 52 78 53
rect -84 36 -82 40
rect -80 36 -77 40
rect -104 4 -102 7
rect -100 4 -98 7
rect -28 49 -24 50
rect -28 44 -24 45
rect 11 44 15 50
rect 40 49 43 50
rect 49 44 52 45
rect 74 44 78 50
rect -28 41 -24 42
rect 11 41 15 42
rect 49 41 52 42
rect 58 36 61 37
rect 74 36 78 42
rect 58 33 61 34
rect 74 33 78 34
rect -8 25 -7 29
rect -4 25 -3 29
rect 34 28 38 29
rect 34 25 38 26
rect 103 25 104 28
rect 106 25 107 28
rect 132 2 133 5
rect 135 2 136 5
<< metal1 >>
rect -87 57 25 60
rect 33 60 60 63
rect 29 57 37 60
rect 40 57 44 60
rect -87 46 -84 57
rect -108 43 -84 46
rect -108 7 -105 43
rect -87 40 -84 43
rect -35 40 -32 57
rect 49 49 52 60
rect 56 57 135 60
rect -24 46 -9 49
rect -35 37 -28 40
rect -77 30 -73 36
rect -77 26 -65 30
rect -77 21 -73 26
rect -68 22 -65 26
rect -12 29 -9 46
rect -68 19 -48 22
rect -68 18 -65 19
rect -88 13 -85 17
rect -42 10 -38 14
rect -3 16 0 25
rect 4 17 7 19
rect 11 17 14 37
rect 40 33 44 45
rect 58 41 61 57
rect 49 33 53 37
rect 38 29 58 33
rect 4 16 22 17
rect -3 14 22 16
rect 34 17 37 21
rect 74 18 78 29
rect 99 29 102 57
rect 108 20 111 25
rect 74 17 90 18
rect 34 15 90 17
rect 108 17 118 20
rect 34 14 78 15
rect -3 13 7 14
rect -42 6 -26 10
rect -3 4 0 13
rect 4 10 7 13
rect -98 -3 -94 3
rect -81 0 -76 4
rect -55 -2 -31 1
rect -98 -4 -86 -3
rect -98 -6 -79 -4
rect -98 -7 -94 -6
rect -90 -7 -79 -6
rect -44 -7 -41 -2
rect -82 -9 -79 -7
rect -107 -27 -104 -11
rect -82 -12 -58 -9
rect -38 -10 -28 -7
rect -88 -27 -85 -14
rect -38 -27 -35 -10
rect -12 -16 -9 0
rect 11 -7 14 14
rect 18 10 21 14
rect 34 11 37 14
rect 74 2 78 14
rect 108 13 111 17
rect 88 6 90 10
rect 38 -1 59 1
rect 34 -2 59 -1
rect 40 -6 43 -2
rect 40 -9 50 -6
rect 40 -15 43 -9
rect -24 -19 -9 -16
rect -107 -30 25 -27
rect 29 -30 36 -27
rect 33 -31 36 -30
rect 39 -31 43 -27
rect 50 -27 54 -19
rect 60 -27 64 -11
rect 99 -27 102 9
rect 128 6 131 57
rect 139 16 149 19
rect 137 -3 140 2
rect 137 -6 145 -3
rect 137 -9 140 -6
rect 128 -27 131 -13
rect 50 -30 131 -27
rect 50 -31 58 -30
rect 33 -34 58 -31
<< metal2 >>
rect 122 16 135 20
rect -88 -10 -85 9
rect 22 6 84 10
<< ntransistor >>
rect -82 17 -80 21
rect -68 -2 -66 1
rect -102 -10 -100 -7
rect 104 10 106 13
rect 34 4 38 6
rect -7 0 -4 4
rect -51 -12 -48 -9
rect 60 -5 63 -3
rect 74 -6 78 -3
rect -28 -14 -24 -12
rect 11 -14 15 -12
rect 51 -14 54 -12
rect 74 -14 78 -12
rect 133 -12 135 -9
rect -28 -22 -24 -20
rect 11 -22 15 -20
rect 40 -22 43 -20
rect 74 -22 78 -20
<< ptransistor >>
rect -28 50 -24 52
rect 11 50 15 52
rect 40 50 43 52
rect 74 50 78 52
rect -82 36 -80 40
rect -102 4 -100 7
rect -28 42 -24 44
rect 11 42 15 44
rect 49 42 52 44
rect 74 42 78 44
rect 58 34 61 36
rect 74 34 78 36
rect -7 25 -4 29
rect 34 26 38 28
rect 104 25 106 28
rect 133 2 135 5
<< polycontact >>
rect -51 15 -47 19
rect -42 14 -38 18
rect -68 5 -64 9
rect -86 0 -81 4
rect -26 6 -22 10
rect 22 14 26 18
rect 90 15 94 19
rect 90 6 94 10
rect -31 -3 -27 1
<< ndcontact >>
rect -88 17 -84 21
rect -77 17 -73 21
rect -76 -2 -71 4
rect -60 -2 -55 3
rect -108 -11 -104 -7
rect -98 -11 -94 -7
rect -58 -12 -53 -7
rect 34 7 38 11
rect 99 9 103 13
rect 107 9 111 13
rect -12 0 -8 4
rect -3 0 1 4
rect 34 -1 38 3
rect 59 -2 63 2
rect 74 -2 78 2
rect -46 -12 -41 -7
rect -28 -11 -24 -7
rect 11 -11 15 -7
rect 50 -10 54 -6
rect 60 -11 64 -7
rect 128 -13 132 -9
rect 136 -13 140 -9
rect -28 -19 -24 -15
rect 39 -19 43 -15
rect 50 -19 54 -15
rect -28 -27 -24 -23
rect 11 -27 15 -23
rect 39 -27 43 -23
rect 74 -27 78 -23
<< pdcontact >>
rect -28 53 -24 57
rect 11 53 15 57
rect 40 53 44 57
rect 74 53 78 57
rect -88 36 -84 40
rect -77 36 -73 40
rect -108 3 -104 7
rect -98 3 -94 7
rect -28 45 -24 49
rect 40 45 44 49
rect 49 45 53 49
rect -28 37 -24 41
rect 11 37 15 41
rect 49 37 53 41
rect 58 37 62 41
rect 34 29 38 33
rect 58 29 62 33
rect 74 29 78 33
rect -12 25 -8 29
rect -3 25 1 29
rect 99 25 103 29
rect 107 25 111 29
rect 34 21 38 25
rect 128 2 132 6
rect 136 2 140 6
<< m2contact >>
rect -88 9 -84 13
rect -89 -14 -85 -10
rect 18 6 22 10
rect 118 16 122 20
rect 84 6 88 10
rect 135 16 139 20
<< psubstratepcontact >>
rect 25 -30 29 -26
<< nsubstratencontact >>
rect 25 57 29 61
<< labels >>
rlabel polysilicon -34 16 -34 16 1 a
rlabel polysilicon -6 16 -6 16 1 c
rlabel metal1 6 59 6 59 5 Vdd
rlabel metal1 2 -29 2 -29 1 Gnd
rlabel polysilicon -81 32 -81 32 1 add
rlabel polysilicon -101 2 -101 2 1 b
rlabel metal1 143 -4 143 -4 7 x
rlabel metal1 148 18 148 18 1 z
<< end >>
