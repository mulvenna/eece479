magic
tech scmos
timestamp 1428795971
<< polysilicon >>
rect 74 139 198 141
rect 74 112 77 139
rect -31 110 77 112
rect -31 16 -28 110
rect 184 17 187 139
rect -94 14 -8 16
rect 184 14 232 17
rect 140 -13 142 -1
rect -94 -15 232 -13
rect -39 -26 196 -24
rect -39 -87 -37 -26
rect -5 -149 -3 -109
rect -94 -499 -16 -496
rect 155 -499 232 -496
rect -94 -508 -17 -505
rect 155 -508 232 -505
rect -94 -545 -17 -543
rect 156 -545 232 -543
rect -19 -714 -17 -697
rect -94 -717 -17 -714
rect 155 -714 157 -697
rect 155 -717 232 -714
<< metal1 >>
rect 174 68 195 69
rect 174 65 196 68
rect 192 -24 196 65
rect -17 -37 -15 -34
rect -11 -37 -9 -34
rect -10 -51 10 -47
rect -87 -131 -82 -53
rect 7 -65 10 -51
rect -60 -72 -45 -68
rect 7 -69 24 -65
rect -62 -73 -45 -72
rect 212 -78 228 -75
rect 208 -131 212 -97
rect -87 -135 212 -131
rect 71 -143 228 -139
rect 53 -389 57 -380
rect 67 -389 71 -381
rect 81 -389 85 -381
rect -94 -400 -17 -396
rect 155 -400 232 -396
rect -94 -409 -17 -405
rect 155 -409 232 -405
rect -94 -419 -17 -415
rect 155 -419 232 -415
rect -94 -429 -17 -425
rect 155 -429 232 -425
rect -94 -439 -17 -435
rect 155 -439 232 -435
rect 82 -456 101 -453
rect 82 -464 85 -456
rect -94 -473 -17 -469
rect 155 -473 232 -469
rect -94 -534 -82 -530
rect -77 -534 39 -530
rect 100 -534 232 -530
rect 75 -743 79 -740
<< metal2 >>
rect -21 -6 -18 13
rect -21 -11 1 -6
rect -55 -51 -14 -47
rect -81 -72 -64 -68
rect -81 -73 -62 -72
rect -81 -530 -77 -73
rect -55 -744 -52 -51
rect -4 -117 0 -11
rect 23 -33 26 -7
rect 21 -84 25 -47
rect -4 -120 2 -117
rect 67 -377 71 -143
rect 149 -148 153 -125
rect 228 -139 232 -78
rect 124 -152 153 -148
rect 85 -381 105 -377
rect 101 -452 105 -381
rect 124 -396 128 -152
rect -55 -747 75 -744
<< polycontact >>
rect 24 -69 28 -65
<< m2contact >>
rect -18 9 -14 13
rect -15 -37 -11 -33
rect 22 -37 26 -33
rect -87 -53 -82 -47
rect -14 -51 -10 -47
rect -64 -72 -60 -68
rect 228 -78 232 -74
rect 21 -88 25 -84
rect -2 -124 2 -120
rect 149 -125 153 -121
rect 67 -143 71 -139
rect 228 -143 232 -139
rect 67 -381 71 -377
rect 81 -381 85 -377
rect 124 -400 128 -396
rect 101 -456 105 -452
rect -82 -535 -77 -530
rect 75 -747 80 -743
use ../cells/reg1  reg1_0
timestamp 1428701549
transform 1 0 35 0 1 37
box -52 -48 141 101
use ../cells/addsub1  addsub1_0
timestamp 1428786523
transform 1 0 63 0 1 -94
box -113 -34 149 63
use dbitlow  dbitlow_0
timestamp 1428705999
transform 1 0 40 0 1 -448
box -57 -292 116 69
<< end >>
