magic
tech scmos
timestamp 1428033508
<< polysilicon >>
rect -8 18 -6 20
rect 7 18 9 20
rect -8 -2 -6 15
rect 7 -2 9 15
rect -8 -7 -6 -5
rect 7 -7 9 -5
<< ndiffusion >>
rect -9 -5 -8 -2
rect -6 -5 7 -2
rect 9 -5 10 -2
<< pdiffusion >>
rect -9 15 -8 18
rect -6 15 -1 18
rect 3 15 7 18
rect 9 15 10 18
<< metal1 >>
rect -13 19 -9 21
rect 10 19 14 21
rect -1 9 3 14
rect -1 6 15 9
rect 10 -1 14 6
rect -13 -7 -9 -5
<< ntransistor >>
rect -8 -5 -6 -2
rect 7 -5 9 -2
<< ptransistor >>
rect -8 15 -6 18
rect 7 15 9 18
<< ndcontact >>
rect -13 -5 -9 -1
rect 10 -5 14 -1
<< pdcontact >>
rect -13 15 -9 19
rect -1 14 3 18
rect 10 15 14 19
<< end >>
