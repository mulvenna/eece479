magic
tech scmos
timestamp 1428795852
<< pwell >>
rect 681 494 717 510
<< nwell >>
rect 681 514 706 536
<< polysilicon >>
rect 689 528 692 536
rect 743 -41 745 -30
rect 752 -41 754 -23
rect 763 -40 765 -16
rect 760 -42 765 -40
rect 768 -42 770 -9
rect 776 -43 778 -34
<< metal1 >>
rect 22 531 678 536
rect 684 530 698 535
rect 703 530 736 535
rect 684 528 688 530
rect 73 524 80 528
rect 236 524 243 528
rect 399 523 406 527
rect 562 523 569 527
rect 736 526 743 530
rect 678 510 693 514
rect 684 499 688 500
rect 684 496 706 499
rect 79 -26 83 0
rect 195 -19 198 0
rect 358 -12 361 3
rect 731 0 780 4
rect 521 -5 524 0
rect 521 -8 766 -5
rect 358 -15 761 -12
rect 195 -22 750 -19
rect 79 -29 741 -26
rect 776 -30 780 0
rect 796 -37 800 24
rect 813 -59 816 -56
<< metal2 >>
rect 812 243 815 332
rect 812 210 815 214
rect 812 162 815 166
rect 741 0 745 4
rect 811 -3 815 0
rect 741 -74 745 -8
<< metal3 >>
rect 739 17 747 19
rect 739 13 741 17
rect 745 13 747 17
rect 739 -4 747 13
rect 739 -8 741 -4
rect 745 -8 747 -4
rect 739 -10 747 -8
<< polycontact >>
rect 80 524 84 528
rect 243 524 247 528
rect 406 523 410 527
rect 569 523 573 527
rect 732 526 736 530
rect 766 -9 770 -5
rect 761 -16 765 -12
rect 750 -23 754 -19
rect 741 -30 745 -26
rect 776 -34 780 -30
<< m2contact >>
rect 741 -78 745 -74
<< m3contact >>
rect 741 13 745 17
rect 741 -8 745 -4
<< nsubstratencontact >>
rect 698 530 703 535
use cvbit  cvbit_0
timestamp 1428795827
transform 1 0 10 0 1 109
box -10 -109 153 422
use cvbit  cvbit_1
timestamp 1428795827
transform 1 0 173 0 1 109
box -10 -109 153 422
use cvbit  cvbit_2
timestamp 1428795827
transform 1 0 336 0 1 109
box -10 -109 153 422
use cvbit  cvbit_3
timestamp 1428795827
transform 1 0 499 0 1 109
box -10 -109 153 422
use ../cells/not  not_0
timestamp 1428691164
transform 1 0 684 0 1 502
box 0 -2 13 26
use cvbit  cvbit_4
timestamp 1428795827
transform 1 0 662 0 1 109
box -10 -109 153 422
use and5  and5_0
timestamp 1428726019
transform 1 0 747 0 1 -81
box -13 0 66 46
<< labels >>
rlabel metal2 813 285 813 285 7 Gnd
rlabel metal2 813 212 813 212 7 clk
rlabel metal2 813 164 813 164 7 Vdd
rlabel metal1 681 512 681 512 1 startb
rlabel polysilicon 690 529 690 529 1 start
rlabel metal1 815 -58 815 -58 7 valid
rlabel metal2 813 -2 813 -2 7 reset
<< end >>
