magic
tech scmos
timestamp 1428796011
<< polysilicon >>
rect 2660 791 2664 802
rect 2710 745 2713 801
rect 2439 458 2442 611
rect 2710 566 2713 743
rect 3853 495 4180 497
rect 2439 454 3783 458
rect 4178 204 4180 495
rect 4092 201 4180 204
<< metal1 >>
rect 402 827 406 1130
rect 729 827 733 1130
rect 1053 827 1057 1130
rect 1380 827 1384 1130
rect 1706 827 1710 1130
rect 2032 827 2036 1130
rect 2358 827 2362 1130
rect 402 824 414 827
rect 729 824 741 827
rect 1053 824 1065 827
rect 1380 824 1392 827
rect 1706 824 1718 827
rect 2032 824 2044 827
rect 2358 824 2370 827
rect 2660 807 2665 1130
rect 2710 806 2715 1129
rect 3836 1128 3842 1129
rect 3749 1127 3842 1128
rect 2764 1123 3842 1127
rect 2764 1120 2774 1123
rect 2764 1075 2772 1120
rect 3836 1061 3842 1123
rect 3841 1055 3842 1061
rect 3756 965 3763 1054
rect 3797 1022 4008 1029
rect 2686 787 2814 791
rect 2740 786 2814 787
rect 2867 788 2925 793
rect 2699 772 2735 776
rect 2719 752 2850 756
rect 2868 749 2873 788
rect 2682 739 2686 748
rect 2868 739 2872 749
rect 2682 734 2872 739
rect 2715 560 2728 561
rect 2710 555 2728 560
rect 2765 504 2772 576
rect 3733 496 3756 499
rect 3752 490 3756 496
rect 3783 460 3788 542
rect 3849 501 3853 542
rect 3888 507 3893 542
rect 3940 516 3945 552
rect 4034 542 4038 1102
rect 3969 529 3973 542
rect 3997 537 4038 542
rect 3969 524 4220 529
rect 3940 513 4200 516
rect 3940 512 3945 513
rect 3888 502 4185 507
rect 3816 486 4225 490
rect 4034 433 4225 437
rect 4034 425 4225 429
rect 4034 417 4225 421
rect 4034 409 4225 413
rect 4034 401 4225 405
rect 4034 393 4225 397
rect 4034 385 4225 389
rect 4034 377 4225 381
rect 4175 341 4201 345
rect 4189 340 4205 341
rect 4209 292 4225 293
rect 4170 288 4221 292
rect 4169 271 4186 275
rect 197 -5 201 3
rect 523 -5 527 3
rect 849 -5 853 2
rect 1175 -5 1179 3
rect 1501 -5 1505 0
rect 1827 -5 1831 1
rect 2153 -5 2157 2
rect 2728 -5 2732 3
rect 2900 -5 2904 4
rect 3072 -5 3076 3
rect 3244 -5 3248 2
rect 3416 -5 3420 10
rect 3588 -5 3592 2
rect 3760 -5 3764 10
rect 3932 -5 3936 10
<< metal2 >>
rect 2734 1102 4029 1106
rect 2734 1101 3820 1102
rect 2734 776 2740 1101
rect 2764 993 2772 1062
rect 3763 1061 3833 1063
rect 3764 1054 3833 1061
rect 3763 1053 3833 1054
rect 4016 1022 4225 1027
rect 2734 775 2735 776
rect 2765 586 2772 993
rect 3763 961 3798 965
rect 2815 717 2820 786
rect 2909 755 2914 764
rect 2857 751 2914 755
rect 2815 713 2915 717
rect 2904 712 2915 713
rect 2734 555 2914 559
rect 3756 486 3812 490
rect 4012 433 4029 437
rect 4012 425 4029 429
rect 4012 417 4029 421
rect 4012 409 4029 413
rect 4012 401 4029 405
rect 4012 393 4029 397
rect 4012 385 4029 389
rect 4012 377 4029 381
rect 4187 275 4190 502
rect 4202 345 4205 512
rect 4222 292 4225 524
<< polycontact >>
rect 2659 802 2665 807
rect 2709 801 2715 806
rect 2710 560 2715 566
rect 3849 495 3853 501
rect 3783 454 3788 460
<< m2contact >>
rect 2764 1062 2773 1075
rect 4029 1102 4038 1108
rect 3756 1054 3764 1061
rect 3833 1054 3841 1061
rect 4008 1022 4016 1029
rect 3756 961 3763 965
rect 3798 961 3802 965
rect 2814 786 2823 791
rect 2735 772 2740 776
rect 2850 751 2857 756
rect 2765 576 2773 586
rect 2728 555 2734 561
rect 3752 486 3756 490
rect 4220 524 4225 529
rect 4200 512 4205 517
rect 4185 502 4190 507
rect 3812 486 3816 490
rect 4029 433 4034 437
rect 4029 425 4034 429
rect 4029 417 4034 421
rect 4029 409 4034 413
rect 4029 401 4034 405
rect 4029 393 4034 397
rect 4029 385 4034 389
rect 4029 377 4034 381
rect 4201 341 4205 345
rect 4221 288 4225 292
rect 4186 271 4190 275
use controller  controller_0
timestamp 1428795880
transform 1 0 2841 0 1 1062
box 73 -588 1184 33
use datapath  datapath_0
timestamp 1428795988
transform 1 0 22 0 1 -38
box -22 38 4164 937
<< labels >>
rlabel metal1 2727 736 2727 736 1 Gnd
rlabel metal1 3934 7 3934 7 1 quotient_0
rlabel metal1 3761 7 3761 7 1 quotient_1
rlabel metal1 3590 -1 3590 -1 1 quotient_2
rlabel metal1 3418 8 3418 8 1 quotient_3
rlabel metal1 3246 -1 3246 -1 1 quotient_4
rlabel metal1 3074 1 3074 1 1 quotient_5
rlabel metal1 2902 1 2902 1 1 quotient_6
rlabel metal1 2730 0 2730 0 1 quotient_7
rlabel metal1 2155 0 2155 0 1 remainder_0
rlabel metal1 1829 -2 1829 -2 1 remainder_1
rlabel metal1 1503 -2 1503 -2 1 remainder_2
rlabel metal1 1177 1 1177 1 1 remainder_3
rlabel metal1 850 -1 850 -1 1 remainder_4
rlabel metal1 525 1 525 1 1 remainder_5
rlabel metal1 199 1 199 1 1 remainder_6
rlabel metal1 2774 736 2774 736 1 Gnd
rlabel metal2 2819 715 2819 715 1 Vdd
rlabel metal1 4219 435 4219 435 1 dividendin_7
rlabel metal1 4218 427 4218 427 1 dividendin_6
rlabel metal1 4218 419 4218 419 1 dividendin_5
rlabel metal1 4218 411 4218 411 1 dividendin_4
rlabel metal1 4217 403 4217 403 1 dividendin_3
rlabel metal1 4217 395 4217 395 1 dividendin_2
rlabel metal1 4217 387 4217 387 1 dividendin_1
rlabel metal1 4217 379 4217 379 1 dividendin_0
rlabel metal1 2360 1125 2360 1125 5 divisorin_0
rlabel metal1 1708 1126 1708 1126 5 divisorin_2
rlabel metal1 2034 1126 2034 1126 5 divisorin_1
rlabel metal1 1382 1125 1382 1125 5 divisorin_3
rlabel metal1 1055 1125 1055 1125 5 divisorin_4
rlabel metal1 731 1126 731 1126 5 divisorin_5
rlabel metal1 404 1127 404 1127 5 divisorin_6
rlabel metal1 2712 1126 2712 1126 5 reset
rlabel metal1 2662 1125 2662 1125 5 clk
rlabel metal2 4219 1024 4219 1024 1 start
rlabel metal1 4215 488 4215 488 1 valid
<< end >>
