magic
tech scmos
timestamp 1428786731
<< pwell >>
rect 38 44 79 58
rect -25 5 18 10
rect 69 5 100 13
rect -25 -8 100 5
rect -73 -9 72 -8
rect -73 -23 1 -9
rect 10 -14 53 -9
rect 13 -67 53 -58
rect -27 -74 53 -67
rect -28 -82 53 -74
rect -28 -87 49 -82
<< nwell >>
rect 32 78 73 81
rect 17 63 73 78
rect 17 38 33 63
rect -32 36 45 38
rect -67 30 45 36
rect -67 20 55 30
rect -67 19 -26 20
rect -75 18 -26 19
rect -75 1 -34 18
rect 14 12 55 20
rect -34 -48 56 -31
rect -34 -62 6 -48
<< polysilicon >>
rect 52 69 55 72
rect 52 63 55 66
rect 37 60 55 63
rect 52 56 55 60
rect 52 38 55 53
rect 52 36 90 38
rect 60 35 90 36
rect 76 12 79 18
rect -49 6 -46 9
rect 88 9 90 35
rect 76 3 79 8
rect -49 -10 -46 3
rect -2 -1 0 3
rect 87 2 90 9
rect -49 -17 -46 -13
rect 45 -22 47 -5
rect 87 -6 90 -2
rect 45 -25 61 -22
rect -3 -36 -2 -32
rect -19 -52 -17 -45
rect -4 -52 -2 -36
rect 43 -41 45 -34
rect 59 -48 61 -25
<< ndiffusion >>
rect 50 53 52 56
rect 55 53 58 56
rect 74 8 76 12
rect 79 8 81 12
rect 85 -2 87 2
rect 90 -2 92 2
rect -51 -13 -49 -10
rect -46 -13 -45 -10
<< pdiffusion >>
rect 50 66 52 69
rect 55 66 58 69
rect -51 3 -49 6
rect -46 3 -45 6
<< metal1 >>
rect 25 76 71 79
rect 25 35 29 76
rect 46 70 49 76
rect 58 62 62 66
rect 58 58 72 62
rect 58 56 62 58
rect 46 49 50 52
rect 37 48 63 49
rect 68 48 72 58
rect 37 45 58 48
rect 62 45 63 48
rect -65 31 -55 35
rect -51 31 -36 35
rect -32 31 56 35
rect -22 29 -18 31
rect 1 29 5 31
rect -70 21 -17 22
rect -70 18 -21 21
rect -61 -3 -58 18
rect 25 20 28 31
rect 48 21 51 31
rect 72 22 76 48
rect 5 15 14 19
rect 72 18 75 22
rect -55 7 -51 10
rect 11 11 14 15
rect 11 7 26 11
rect 53 8 70 11
rect 85 8 120 11
rect -61 -6 -53 -3
rect -45 -4 -41 3
rect -28 1 -18 4
rect 68 -1 81 2
rect -45 -5 -20 -4
rect -45 -8 -21 -5
rect -45 -10 -41 -8
rect -69 -20 -64 -17
rect -55 -17 -51 -14
rect -60 -20 -10 -17
rect -59 -56 -55 -20
rect -36 -24 -31 -23
rect -2 -24 1 -5
rect 25 -9 29 -5
rect 68 -9 71 -1
rect 96 -1 99 8
rect 102 6 120 8
rect 25 -13 28 -9
rect 25 -17 29 -13
rect 9 -20 29 -17
rect -37 -28 1 -24
rect -36 -64 -31 -28
rect 102 -30 105 6
rect -16 -35 -7 -32
rect 46 -34 106 -30
rect 58 -35 106 -34
rect 0 -40 6 -37
rect 10 -40 50 -37
rect 0 -47 3 -40
rect 23 -41 27 -40
rect 46 -41 50 -40
rect -24 -50 3 -47
rect -24 -53 -20 -50
rect -1 -53 3 -50
rect 12 -55 24 -52
rect 51 -55 84 -52
rect 12 -63 16 -55
rect -72 -68 -23 -64
rect 4 -66 16 -63
rect -24 -80 -20 -79
rect 23 -80 27 -68
rect -28 -82 17 -80
rect -55 -84 17 -82
rect 21 -84 48 -80
rect -55 -85 48 -84
<< metal2 >>
rect 15 45 33 48
rect -70 -47 -66 31
rect -55 14 -51 31
rect -32 -13 -28 1
rect -20 -31 -15 -11
rect 15 -13 19 45
rect 33 -13 67 -9
rect -6 -20 5 -17
rect -70 -51 -28 -47
rect -59 -81 -56 -60
<< ntransistor >>
rect 52 53 55 56
rect 76 8 79 12
rect 87 -2 90 2
rect -49 -13 -46 -10
<< ptransistor >>
rect 52 66 55 69
rect -49 3 -46 6
<< polycontact >>
rect 72 48 76 52
rect -21 17 -17 21
rect 75 18 79 22
rect 26 7 30 11
rect -53 -6 -49 -2
rect -3 -5 1 -1
rect -7 -36 -3 -32
rect 42 -34 46 -30
rect 24 -55 28 -51
rect 57 -52 61 -48
rect -23 -68 -19 -64
<< ndcontact >>
rect 46 52 50 56
rect 58 52 62 56
rect 70 8 74 12
rect 81 8 85 12
rect 81 -2 85 2
rect 92 -2 96 2
rect -55 -14 -51 -10
rect -45 -14 -41 -10
<< pdcontact >>
rect 46 66 50 70
rect 58 66 62 70
rect -55 3 -51 7
rect -45 3 -41 7
<< m2contact >>
rect 33 45 37 49
rect -70 31 -65 35
rect -55 31 -51 35
rect -55 10 -51 14
rect -32 1 -28 5
rect -21 -11 -16 -5
rect -32 -17 -28 -13
rect -10 -20 -6 -16
rect 28 -13 33 -9
rect 67 -13 72 -9
rect 5 -20 9 -16
rect 15 -17 19 -13
rect -59 -60 -55 -56
rect -20 -35 -16 -31
rect -28 -51 -24 -47
rect -59 -85 -55 -81
<< psubstratepcontact >>
rect 58 44 62 48
rect -64 -20 -60 -16
rect 17 -84 21 -80
<< nsubstratencontact >>
rect -36 31 -32 35
rect 6 -40 10 -36
use nand  nand_0
timestamp 1428033508
transform 1 0 -9 0 1 10
box -13 -7 15 21
use nand  nand_1
timestamp 1428033508
transform 1 0 38 0 1 2
box -13 -7 15 21
use nand  nand_2
timestamp 1428033508
transform 1 0 -11 0 1 -72
box -13 -7 15 21
use nand  nand_3
timestamp 1428033508
transform 1 0 36 0 1 -61
box -13 -7 15 21
<< labels >>
rlabel metal1 -71 -66 -71 -66 3 clk
rlabel polysilicon 38 62 38 62 1 reset
rlabel metal1 -68 20 -68 20 3 d
rlabel metal1 104 10 104 10 7 q
rlabel metal1 -20 33 -20 33 1 Vdd
rlabel metal1 -36 -83 -36 -83 1 Gnd
<< end >>
