magic
tech scmos
timestamp 1428530478
<< pwell >>
rect -25 -19 25 0
<< nwell >>
rect -25 5 25 24
<< polysilicon >>
rect -20 16 -16 24
rect -3 16 1 24
rect 11 13 18 16
rect 23 13 25 16
rect -20 0 -16 12
rect -20 -7 -16 -4
rect -3 11 1 12
rect -3 -7 1 7
rect 11 5 15 13
rect 11 -8 15 0
rect 11 -11 18 -8
rect 23 -11 25 -8
rect -20 -19 -16 -11
rect -3 -19 1 -11
<< ndiffusion >>
rect -21 -11 -20 -7
rect -16 -11 -11 -7
rect -7 -11 -3 -7
rect 1 -11 4 -7
rect 18 -8 23 -7
rect 18 -15 23 -11
<< pdiffusion >>
rect 18 16 23 20
rect -21 12 -20 16
rect -16 12 -3 16
rect 1 12 4 16
rect 18 12 23 13
<< metal1 >>
rect -25 20 9 24
rect 13 20 18 24
rect 23 20 25 24
rect -25 16 -21 20
rect -18 9 -3 11
rect -25 7 -3 9
rect -25 5 -14 7
rect 4 5 8 12
rect 18 5 23 8
rect 4 4 11 5
rect -11 0 11 4
rect 18 0 25 5
rect -25 -4 -20 0
rect -11 -7 -7 0
rect 18 -3 23 0
rect -25 -15 -21 -11
rect 4 -15 8 -11
rect -25 -19 9 -15
rect 13 -19 18 -15
rect 23 -19 25 -15
<< ntransistor >>
rect -20 -11 -16 -7
rect -3 -11 1 -7
rect 18 -11 23 -8
<< ptransistor >>
rect -20 12 -16 16
rect -3 12 1 16
rect 18 13 23 16
<< polycontact >>
rect -20 -4 -16 0
rect -3 7 1 11
rect 11 0 15 5
<< ndcontact >>
rect -25 -11 -21 -7
rect -11 -11 -7 -7
rect 4 -11 8 -7
rect 18 -7 23 -3
rect 18 -19 23 -15
<< pdcontact >>
rect 18 20 23 24
rect -25 12 -21 16
rect 4 12 8 16
rect 18 8 23 12
<< psubstratepcontact >>
rect 9 -19 13 -15
<< nsubstratencontact >>
rect 9 20 13 24
<< labels >>
rlabel metal1 24 2 24 2 7 z
rlabel polysilicon -2 5 -2 6 5 b
rlabel polysilicon -17 3 -17 3 5 a
rlabel metal1 -24 23 -24 23 4 Vdd
rlabel metal1 -24 -18 -24 -18 2 Gnd
<< end >>
