magic
tech scmos
timestamp 1428691952
<< polysilicon >>
rect 1 7 3 9
rect 1 -1 3 1
rect 1 -9 3 -7
rect 1 -14 3 -12
<< ndiffusion >>
rect 0 -12 1 -9
rect 3 -12 4 -9
<< pdiffusion >>
rect 0 1 1 7
rect 3 1 4 7
<< metal1 >>
rect -4 -2 0 1
rect -7 -6 0 -2
rect -4 -9 0 -6
rect 4 -2 8 1
rect 4 -6 11 -2
rect 4 -9 8 -6
<< ntransistor >>
rect 1 -12 3 -9
<< ptransistor >>
rect 1 1 3 7
<< ndcontact >>
rect -4 -13 0 -9
rect 4 -13 8 -9
<< pdcontact >>
rect -4 1 0 7
rect 4 1 8 7
<< end >>
