magic
tech scmos
timestamp 1428029823
<< pwell >>
rect -25 -19 25 1
<< nwell >>
rect -25 4 25 24
<< polysilicon >>
rect -20 16 -16 24
rect -3 16 1 24
rect 11 13 18 16
rect 23 13 25 16
rect -20 9 -16 12
rect -20 -7 -16 5
rect -3 -2 1 12
rect -3 -7 1 -6
rect 11 5 15 13
rect 11 -8 15 0
rect 11 -11 18 -8
rect 23 -11 25 -8
rect -20 -19 -16 -11
rect -3 -19 1 -11
<< ndiffusion >>
rect -21 -11 -20 -7
rect -16 -11 -3 -7
rect 1 -11 4 -7
rect 18 -8 23 -7
rect 18 -15 23 -11
<< pdiffusion >>
rect 18 16 23 20
rect -21 12 -20 16
rect -16 12 -11 16
rect -7 12 -3 16
rect 1 12 4 16
rect 18 12 23 13
<< metal1 >>
rect -25 20 9 24
rect 13 20 18 24
rect 23 20 25 24
rect -25 16 -21 20
rect 4 16 8 20
rect -25 5 -20 9
rect -11 5 -7 12
rect 18 5 23 8
rect -11 1 11 5
rect 4 0 11 1
rect 18 0 25 5
rect -25 -2 -14 0
rect -25 -4 -3 -2
rect -18 -6 -3 -4
rect 4 -7 8 0
rect 18 -3 23 0
rect -25 -15 -21 -11
rect -25 -19 9 -15
rect 13 -19 18 -15
rect 23 -19 25 -15
<< ntransistor >>
rect -20 -11 -16 -7
rect -3 -11 1 -7
rect 18 -11 23 -8
<< ptransistor >>
rect -20 12 -16 16
rect -3 12 1 16
rect 18 13 23 16
<< polycontact >>
rect -20 5 -16 9
rect -3 -6 1 -2
rect 11 0 15 5
<< ndcontact >>
rect -25 -11 -21 -7
rect 4 -11 8 -7
rect 18 -7 23 -3
rect 18 -19 23 -15
<< pdcontact >>
rect 18 20 23 24
rect -25 12 -21 16
rect -11 12 -7 16
rect 4 12 8 16
rect 18 8 23 12
<< psubstratepcontact >>
rect 9 -19 13 -15
<< nsubstratencontact >>
rect 9 20 13 24
<< labels >>
rlabel metal1 24 3 24 3 7 z
rlabel metal1 -23 22 -23 22 4 Vdd
rlabel metal1 -23 -17 -23 -17 2 Gnd
rlabel polysilicon -2 -1 -2 0 1 b
rlabel polysilicon -17 2 -17 2 1 a
<< end >>
