magic
tech scmos
timestamp 1428795880
<< polysilicon >>
rect 762 29 812 33
rect 907 -231 921 -229
rect 1137 -244 1141 -243
rect 1010 -306 1085 -302
rect 888 -368 920 -366
<< metal1 >>
rect 816 29 956 33
rect 936 -176 940 -71
rect 952 -85 956 29
rect 956 -89 967 -85
rect 961 -100 966 -95
rect 1083 -129 1087 -128
rect 1083 -131 1089 -129
rect 1083 -132 1085 -131
rect 1117 -132 1121 -128
rect 944 -202 948 -147
rect 988 -217 991 -194
rect 1014 -223 1019 -171
rect 903 -293 907 -233
rect 1057 -234 1060 -180
rect 1085 -214 1089 -180
rect 1148 -190 1152 -147
rect 1137 -238 1138 -234
rect 1137 -239 1141 -238
rect 944 -256 948 -244
rect 970 -256 974 -244
rect 968 -291 970 -287
rect 967 -292 971 -291
rect 884 -462 888 -370
rect 923 -459 927 -388
rect 975 -459 979 -398
rect 987 -427 991 -400
rect 1035 -435 1038 -378
rect 1052 -431 1056 -430
rect 1061 -451 1065 -294
rect 1118 -368 1122 -356
rect 1118 -426 1122 -398
rect 1176 -431 1180 -404
rect 942 -520 947 -516
rect 1008 -520 1012 -516
rect 1047 -520 1052 -516
rect 1099 -520 1104 -516
rect 1128 -520 1133 -516
rect 1156 -520 1161 -516
rect 889 -566 892 -563
<< metal2 >>
rect 940 -71 1036 -67
rect 870 -80 966 -76
rect 1032 -77 1036 -71
rect 1148 -95 1152 -87
rect 1027 -104 1050 -100
rect 948 -147 966 -143
rect 964 -156 966 -152
rect 1085 -176 1089 -135
rect 940 -180 1056 -176
rect 992 -194 1148 -190
rect 885 -212 923 -209
rect 944 -240 948 -206
rect 970 -206 1151 -202
rect 970 -240 974 -206
rect 1117 -218 1121 -215
rect 885 -297 903 -293
rect 944 -439 948 -260
rect 970 -287 974 -260
rect 1057 -294 1061 -238
rect 1104 -351 1108 -227
rect 1147 -234 1151 -206
rect 1142 -238 1151 -234
rect 1104 -355 1118 -351
rect 1057 -363 1079 -359
rect 1118 -394 1122 -372
rect 1104 -400 1108 -399
rect 1172 -404 1176 -400
rect 1021 -427 1025 -426
rect 991 -431 1021 -427
rect 1056 -430 1118 -426
<< metal3 >>
rect 1102 -83 1154 -81
rect 1102 -87 1148 -83
rect 1152 -87 1154 -83
rect 1102 -89 1154 -87
rect 1020 -100 1029 -99
rect 1020 -104 1023 -100
rect 1027 -104 1029 -100
rect 1020 -105 1029 -104
rect 959 -152 965 -151
rect 959 -156 960 -152
rect 964 -156 965 -152
rect 959 -443 965 -156
rect 1020 -422 1026 -105
rect 1102 -400 1110 -89
rect 1102 -404 1104 -400
rect 1108 -404 1110 -400
rect 1102 -407 1110 -404
rect 1020 -426 1021 -422
rect 1025 -426 1026 -422
rect 1020 -427 1026 -426
rect 959 -447 960 -443
rect 964 -447 965 -443
rect 959 -448 965 -447
<< polycontact >>
rect 812 29 816 33
rect 903 -233 907 -229
rect 1137 -243 1141 -239
rect 967 -296 971 -292
rect 884 -370 888 -366
<< m2contact >>
rect 936 -71 940 -67
rect 866 -80 870 -76
rect 966 -80 970 -76
rect 952 -89 956 -85
rect 1148 -99 1152 -95
rect 1085 -135 1089 -131
rect 936 -180 940 -176
rect 944 -147 948 -143
rect 966 -147 970 -143
rect 966 -156 970 -152
rect 944 -206 948 -202
rect 988 -194 992 -190
rect 923 -212 927 -208
rect 1056 -180 1060 -176
rect 1085 -180 1089 -176
rect 1148 -194 1152 -190
rect 1085 -218 1089 -214
rect 1104 -227 1108 -223
rect 1057 -238 1061 -234
rect 1138 -238 1142 -234
rect 944 -244 948 -240
rect 944 -260 948 -256
rect 970 -244 974 -240
rect 970 -260 974 -256
rect 970 -291 974 -287
rect 903 -297 907 -293
rect 1061 -294 1065 -290
rect 1053 -363 1057 -359
rect 975 -398 979 -394
rect 987 -431 991 -427
rect 1021 -431 1025 -427
rect 1052 -430 1056 -426
rect 1035 -439 1039 -435
rect 1118 -356 1122 -352
rect 1118 -372 1122 -368
rect 1104 -399 1108 -395
rect 1118 -398 1122 -394
rect 1168 -404 1172 -400
rect 1176 -404 1180 -400
rect 1118 -430 1122 -426
rect 1061 -455 1065 -451
<< m3contact >>
rect 1148 -87 1152 -83
rect 1023 -104 1027 -100
rect 960 -156 964 -152
rect 1104 -404 1108 -400
rect 1021 -426 1025 -422
rect 960 -447 964 -443
use cvalid  cvalid_0
timestamp 1428795852
transform 1 0 73 0 1 -507
box 0 -81 816 536
use cnext  cnext_0
timestamp 1428536589
transform 1 0 996 0 1 -174
box -30 3 152 98
use ../cells/reg1  reg1_0
timestamp 1428701549
transform 0 1 959 -1 0 -261
box -52 -48 141 101
use ../cells/reg1  reg1_1
timestamp 1428701549
transform 0 -1 1136 1 0 -351
box -52 -48 141 101
use coutput  coutput_0
timestamp 1428541776
transform 0 1 977 -1 0 -459
box -28 -62 57 203
<< labels >>
rlabel m2contact 989 -429 989 -429 3 c0
rlabel m2contact 1037 -437 1037 -436 3 c0b
rlabel m2contact 1063 -453 1063 -453 3 c1b
rlabel m2contact 1054 -428 1054 -428 3 c1
rlabel metal1 1010 -518 1010 -518 1 shift
rlabel metal1 945 -518 945 -518 1 add
rlabel metal1 1050 -518 1050 -518 1 inbit
rlabel metal1 1102 -519 1102 -519 1 sel1
rlabel metal1 1131 -518 1131 -518 1 sel2
rlabel metal1 1159 -518 1159 -518 1 load
rlabel polysilicon 1048 -304 1048 -304 3 clk
rlabel metal3 1106 -180 1106 -180 3 n1
rlabel m2contact 1150 -192 1150 -192 3 n0
rlabel metal1 962 -97 962 -97 3 sign
rlabel metal2 1148 -204 1148 -204 3 reset
rlabel metal1 1178 -417 1178 -416 3 Gnd
rlabel metal1 925 -415 925 -415 3 Vdd
rlabel metal1 890 -565 890 -565 1 valid
rlabel metal1 954 31 954 31 5 start
<< end >>
