magic
tech scmos
timestamp 1428459501
<< pwell >>
rect -36 -6 25 50
<< nwell >>
rect -36 -22 25 -6
<< polysilicon >>
rect -22 36 -19 45
rect -3 43 1 53
rect -24 32 -19 36
rect 2 28 4 31
rect 8 28 19 31
rect -16 25 -12 28
rect -8 25 -6 28
rect -36 13 12 16
rect 16 13 25 16
rect -36 4 -3 7
rect 1 4 25 7
rect -20 -11 -17 -6
rect 5 -11 8 -8
rect -20 -17 -17 -15
rect 5 -17 8 -15
<< ndiffusion >>
rect 4 31 8 32
rect -12 28 -8 29
rect 4 27 8 28
rect -12 24 -8 25
rect 12 16 16 17
rect 12 12 16 13
rect -3 7 1 8
rect -3 3 1 4
<< pdiffusion >>
rect -21 -15 -20 -11
rect -17 -15 -16 -11
rect 4 -15 5 -11
rect 8 -15 9 -11
<< metal1 >>
rect -36 46 -17 50
rect -13 46 21 50
rect -36 39 -3 43
rect -13 33 -8 36
rect -13 32 -12 33
rect -28 24 -24 32
rect -32 20 -24 24
rect -32 -11 -28 20
rect -20 3 -17 24
rect -12 12 -8 20
rect -3 12 1 39
rect 4 36 8 46
rect 12 39 25 43
rect 4 22 8 23
rect 12 21 16 39
rect 12 3 16 8
rect -20 -1 -3 3
rect 1 -1 16 3
rect -20 -2 -17 -1
rect 19 -4 23 28
rect -8 -8 5 -4
rect 9 -8 23 -4
rect -12 -15 -9 -8
rect 13 -15 19 -11
rect -25 -18 -21 -15
rect 0 -18 4 -15
rect -36 -22 -32 -18
rect -28 -22 21 -18
<< metal2 >>
rect -17 36 -13 46
rect -12 -4 -8 8
rect 4 2 8 18
rect 4 -2 23 2
rect 19 -11 23 -2
rect -32 -18 -28 -15
rect 13 -15 19 -11
rect 13 -21 17 -15
rect 0 -25 17 -21
<< ntransistor >>
rect 4 28 8 31
rect -12 25 -8 28
rect 12 13 16 16
rect -3 4 1 7
<< ptransistor >>
rect -20 -15 -17 -11
rect 5 -15 8 -11
<< polycontact >>
rect -3 53 1 57
rect -3 39 1 43
rect -28 32 -24 36
rect 19 28 23 32
rect -20 24 -16 28
rect -21 -6 -17 -2
rect 5 -8 9 -4
<< ndcontact >>
rect -12 29 -8 33
rect 4 32 8 36
rect -12 20 -8 24
rect 4 23 8 27
rect 12 17 16 21
rect -3 8 1 12
rect 12 8 16 12
rect -3 -1 1 3
<< pdcontact >>
rect -25 -15 -21 -11
rect -16 -15 -12 -11
rect 0 -15 4 -11
rect 9 -15 13 -11
<< m2contact >>
rect -17 46 -13 50
rect -17 32 -13 36
rect -12 8 -8 12
rect 4 18 8 22
rect -12 -8 -8 -4
rect -32 -15 -28 -11
rect 19 -15 23 -11
rect -32 -22 -28 -18
rect 0 -29 4 -25
<< psubstratepcontact >>
rect 21 46 25 50
<< nsubstratencontact >>
rect 21 -22 25 -18
<< labels >>
rlabel polysilicon 24 6 24 6 7 shiftb
rlabel polysilicon 24 15 24 15 7 shift
rlabel nsubstratencontact 24 -19 24 -19 8 Vdd
rlabel m2contact 2 -27 2 -27 1 out
rlabel psubstratepcontact 23 48 23 48 7 Gnd
rlabel metal1 24 41 24 41 7 inbit
rlabel polycontact -1 55 -1 55 5 in
<< end >>
