magic
tech scmos
timestamp 1428690772
<< polysilicon >>
rect -8 23 -6 25
rect 7 23 9 25
rect -8 -1 -6 15
rect 7 -1 9 15
rect -8 -7 -6 -5
rect 7 -7 9 -5
<< ndiffusion >>
rect -9 -5 -8 -1
rect -6 -5 -1 -1
rect 3 -5 7 -1
rect 9 -5 10 -1
<< pdiffusion >>
rect -9 15 -8 23
rect -6 15 7 23
rect 9 15 10 23
<< metal1 >>
rect -13 23 -9 25
rect 10 8 14 15
rect -1 5 15 8
rect -1 -1 3 5
rect -13 -7 -9 -5
rect 10 -7 14 -5
<< ntransistor >>
rect -8 -5 -6 -1
rect 7 -5 9 -1
<< ptransistor >>
rect -8 15 -6 23
rect 7 15 9 23
<< ndcontact >>
rect -13 -5 -9 -1
rect -1 -5 3 -1
rect 10 -5 14 -1
<< pdcontact >>
rect -13 15 -9 23
rect 10 15 14 23
<< end >>
